program test();

  environment env;
  
  initial
    begin
      
      env = new();
      
      env.run();
    end
  
endprogram
  
  
