interface inter_face(input logic clk);
  logic in;
  logic Rise_Detect, Fall_Detect;
  
endinterface
