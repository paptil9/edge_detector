
  `include "transaction.sv"

  `include "interface.sv"

  `include "d_config.sv"

  `include"generator.sv"
  `include"driver.sv"
  `include"pmonitor.sv"
  `include"scoreboard.sv"
  `include "environment.sv"
  `include "test.sv"
  `include "checkerflag.sv"

